// Miren Bamforth | A Motion-Tracking DMX512 Controller
// 6.111 Final Project | Fall 2014
// This code was modified from code on the 6.111 website.

// A high level block which contains everything in the motion
// tracking block to help keep labkit.v cleaner.
module tracking_block(input reset,
								input clk
			);


endmodule
