`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:07:45 11/24/2014 
// Design Name: 
// Module Name:    arctan_lut 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module arctan_lut(
    input clk,
    input reset,
    input [10:0] in,
    output [7:0] out
    );


endmodule
