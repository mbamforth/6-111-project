// Miren Bamforth | A Motion-Tracking DMX512 Controller
// 6.111 Final Project | Fall 2014
// This code was modified from code on the 6.111 website.

//
// File:   zbt_6111.v
// Date:   27-Nov-05
// Author: I. Chuang <ichuang@mit.edu>
//
// Simple ZBT driver for the MIT 6.111 labkit, which does not hide the
// pipeline delays of the ZBT from the user.  The ZBT memories have
// two cycle latencies on read and write, and also need extra-long data hold
// times around the clock positive edge to work reliably.
//

/////////////////////////////////////////////////////////////////////////////
// Ike's simple ZBT RAM driver for the MIT 6.111 labkit
//
// Data for writes can be presented and clocked in immediately; the actual
// writing to RAM will happen two cycles later.
//
// Read requests are processed immediately, but the read data is not available
// until two cycles after the intial request.
//
// A clock enable signal is provided; it enables the RAM clock when high.

module zbt_6111(clk, cen, we, addr, write_data, frame_enable, read_data,
		  ram_clk, ram_we_b, ram_address, ram_data, ram_cen_b);

   input clk;			// system clock
   input cen;			// clock enable for gating ZBT cycles
   input we;			// write enable (active HIGH)
   input [18:0] addr;		// memory address
   input [35:0] write_data;	// data to write
	input frame_enable; // we write every nth frame because of this
   output [35:0] read_data;	// data read from memory
   output 	 ram_clk;	// physical line to ram clock
   output 	 ram_we_b;	// physical line to ram we_b
   output [18:0] ram_address;	// physical line to ram address
   inout [35:0]  ram_data;	// physical line to ram data
   output 	 ram_cen_b;	// physical line to ram clock enable

   // clock enable (should be synchronous and one cycle high at a time)
   wire 	 ram_cen_b = ~cen;

   // create delayed ram_we signal: note the delay is by two cycles!
   // ie we present the data to be written two cycles after we is raised 
   // this means the bus is tri-stated two cycles after we is raised.

   reg [1:0]   we_delay;

   always @(posedge clk)
     we_delay <= cen ? {we_delay[0],we} : we_delay;
   
   // create two-stage pipeline for write data

   reg [35:0]  write_data_old1;
   reg [35:0]  write_data_old2;
   always @(posedge clk)
     if (cen)
       {write_data_old2, write_data_old1} <= {write_data_old1, write_data};

   // wire to ZBT RAM signals
   assign      ram_we_b = ~(we && frame_enable);
	//assign      ram_we_b = ~(we);
	assign      ram_clk = 1'b0;  // gph 2011-Nov-10
	                              // set to zero as place holder
											
//   assign      ram_clk = ~clk;     // RAM is not happy with our data hold
                                   // times if its clk edges equal FPGA's
                                   // so we clock it on the falling edges
                                   // and thus let data stabilize longer
   assign      ram_address = addr;
   
   assign      ram_data = we_delay[1] ? write_data_old2 : {36{1'bZ}};
   assign      read_data = ram_data;

endmodule // zbt_6111

